`define SONG_WIDTH 7
`define NOTE_WIDTH 6
`define DURATION_WIDTH 6
`define METADATA_WIDTH 3


`define SWIDTH 4
`define IDLE   4'b0000
`define LOAD   4'b0001
`define DELAY  4'b0010
`define NOTE1  4'b0011
`define NOTE2  4'b0100
`define NOTE3  4'b0101
`define NOTE4  4'b0110
`define PLAY   4'b0111
`define WAIT   4'b1000

module song_reader(
   input clk,
   input reset,
   input play,
   input [1:0] song,
   input note_done,
   output wire song_done,
   output wire [5:0] note1,
   output wire [5:0] note2, //new additional
   output wire [5:0] note3, //new additional
   output wire [5:0] note4, //new additional
   output wire [5:0] duration, 
   output wire new_note,  
   output wire [1:0] num_notes, //new output
   output wire [2:0] metadata1, //for harmonics
   output wire [2:0] metadata2, //new additional
   output wire [2:0] metadata3, //new additional
   output wire [2:0] metadata4 //new additional
);

    // Declaring wires
    wire [`SONG_WIDTH - 1:0] curr_songaddr, next_songaddr; 
    wire [`SONG_WIDTH + 1:0] rom_addr = {song, curr_songaddr};
    wire [`NOTE_WIDTH + `DURATION_WIDTH + `METADATA_WIDTH:0] note_duration_metadata;

    wire [`SWIDTH-1:0] state;
    reg  [`SWIDTH-1:0] next;


    // ROM for addressing the song
    song_rom rom(.clk(clk), .addr(rom_addr), .dout(note_duration_metadata));


    // Case statements for FSM
    always @(*) begin
        case (state)
            `IDLE:      next = play ? `LOAD : `IDLE; 
            `LOAD:      next = play ? `DELAY : `IDLE; 
            `DELAY:     next = play ? `NOTE1 : `IDLE; 
            `NOTE1:     next = play ? (trigger ? `PLAY : `NOTE2) : `IDLE; 
            `NOTE2:     next = play ? (trigger ? `PLAY : `NOTE3) : `IDLE;
            `NOTE3:     next = play ? (trigger ? `PLAY : `NOTE4) : `IDLE;
            `NOTE4:     next = play ? `PLAY : `IDLE;
            `PLAY:      next = play ? `WAIT : `IDLE;
            `WAIT:      next = note_done ? `IDLE : `WAIT;
            default:    next = `IDLE;
        endcase
    end

    wire trigger;       // For identifying when we should pass time
    wire overflow;      // For identifying when we reach the end of a song
    assign {overflow, next_songaddr} =
       (state == `LOAD || state == `DELAY || state == `NOTE1 || state == `NOTE2) ? {1'b0, curr_songaddr} + 1
                                     : {1'b0, curr_songaddr};

    // To alert notes player that new notes have been added
    assign new_note = (state == `PLAY); 

    wire [5:0] next_duration;
    wire [2:0] metadata;

    assign trigger = note_duration_metadata[15];
    assign note = note_duration_metadata[14:9];
    assign next_duration = note_duration_metadata[8:3];
    assign metadata = note_duration_metadata[2:0];
    assign song_done = overflow;


    // Flip flop for address
    dffre #(`SONG_WIDTH) note_counter (
       .clk(clk),
       .r(reset),
       .en(state <= `NOTE2 && !trigger),
       .d(next_songaddr),
       .q(curr_songaddr)
    );


    // Flip flop for FSM state
    dffr #(`SWIDTH) fsm (
       .clk(clk),
       .r(reset),
       .d(next),
       .q(state)
    );


    // Case statement for number of notes based on state
    reg [1:0] next_num_notes;
    always @(*) begin
        case(state)
            `NOTE1: next_num_notes = 2'b00;
            `NOTE2: next_num_notes = 2'b01;
            `NOTE3: next_num_notes = 2'b10;
            `NOTE4: next_num_notes = 2'b11;
            default: next_num_notes = 2'b00;
        endcase
    end


    // Flip flop for number of notes
    dffre #(2) num_notes_ff (
        .clk(clk),
        .r(reset),
        .en(state < `PLAY),
        .d(next_num_notes),
        .q(num_notes)
    );


    wire [5:0] note;

    // Flip flops for seperate notes
    dffre #(`NOTE_WIDTH + `METADATA_WIDTH) note1_FF(
        .clk(clk), .r(reset || state == `IDLE),
        .en(state == `DELAY), 
        .d({note, metadata}), .q({note1, metadata1})
    );

    dffre #(`NOTE_WIDTH + `METADATA_WIDTH) note2_FF(
        .clk(clk), .r(reset || state == `IDLE),
        .en(state == `NOTE1), 
        .d({note, metadata}), .q({note2, metadata2})
    );

    dffre #(`NOTE_WIDTH + `METADATA_WIDTH) note3_FF(
        .clk(clk), .r(reset || state == `IDLE),
        .en(state == `NOTE2), 
        .d({note, metadata}), .q({note3, metadata3})
    );

    dffre #(`NOTE_WIDTH + `METADATA_WIDTH) note4_FF(
        .clk(clk), .r(reset || state == `IDLE),
        .en(state == `NOTE3), 
        .d({note, metadata}), .q({note4, metadata4})
    );


    // Flip flop for metadata
    // NOTE: we made the assumption that the song rom has chords that have the same metadata and duration
    // Add new_note
    dffre #(`DURATION_WIDTH) metadata_duration_FF(
        .clk(clk), .r(reset || state == `IDLE),
        .en(state == `DELAY),
        .d({next_duration}), .q({duration})
    );

endmodule
